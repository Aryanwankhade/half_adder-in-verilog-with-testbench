`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 28.01.2026 23:48:47
// Design Name: 
// Module Name: full_adders
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module full_adders(a,b,c,sum,carry);
input a,b,c;
output sum ,carry;
assign sum=a^b^c;
assign carry = a&b| b&c | a&c;
endmodule
